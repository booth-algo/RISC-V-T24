module hazard_unit (
    input rst,
);

    // Data hazard

    // Control hazard

    // Stall control

    // Flush control



endmodule
