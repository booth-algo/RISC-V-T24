module controlunit #(
    parameter 
) (
   
);
    
endmodule

// Control Unit is not clocked and decodes the instruction to provide control signals to various modules