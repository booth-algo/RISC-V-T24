module hazard_unit (
    input logic rst,
    input logic [1:0] forwardAE,
    input logic [1:0] forwardBE
    output logic [1:0] forwardAE_out

);

    // Data hazard
    always_comb begin

    end

    // Control hazard

    // Stall control

    // Flush control



endmodule
