module regfile #(
    parameter WIDTH = 32
) (
    input logic     rs1,
    input logic     rs2,
    input logic     rd,
    input logic     RegWrite,
    input logic     ALUout,
    input logic     clk,
    output logic    ALUop1,
    output logic    regOp2
);


    
endmodule